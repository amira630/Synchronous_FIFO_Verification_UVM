package fifo_transactions_pkg;

    // Standard UVM import & include:
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import shared_pkg::*;
    
    // Includes:
    `include "fifo_config.svh"
    `include "fifo_seq_item.svh"

endpackage