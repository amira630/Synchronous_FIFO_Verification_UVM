//////////////////////////////////////////////////////////////////////////////////////////////////////
// Author: Amira Atef
// Course: Digital Verification using SV & UVM
// Date: 04-07-2025
// Description: Package containing shared types and variables for the FIFO verification environment
//////////////////////////////////////////////////////////////////////////////////////////////////////

package shared_pkg;
    bit test_finished; // Flag to indicate if the test is finished

    ////////////////////////////////////////////////////////
    ////////////////////// Counters ////////////////////////
    ////////////////////////////////////////////////////////

    int correct_count, error_count;

    /////////////////////////////////////////////////////////
    ///////////////////// Parameters ////////////////////////
    /////////////////////////////////////////////////////////

    parameter int FIFO_WIDTH = 16; // Width of the FIFO data bus
    parameter int FIFO_DEPTH = 8; // Depth of the FIFO
endpackage